 module enemies(
    input wire pclk,                                  // Peripheral Clock
    input wire rst,                                   // Synchrous reset


    output wire [3:0] level,
  );

  endmodule